module fpu_add_sub();

	input [31:0]floating1;
	input [31:0]floating2;
	
	output [31:0]floating_result;
	
	wire 
	
	
endmodule 