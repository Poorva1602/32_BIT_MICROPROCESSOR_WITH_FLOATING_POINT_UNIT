module control();

	input 
	
	output 


endmodule